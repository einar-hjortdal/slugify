module slugify

const substitutions_no = {
	'&': 'og'
	'@': 'at'
	'æ': 'ae'
	'ø': 'oe'
	'å': 'aa'
	'Æ': 'Ae'
	'Ø': 'Oe'
	'Å': 'Aa'
}
