module slugify

// `en` should always be the first in the map.
const language_to_substitutions = {
	'en': substitutions_en
	'fa': substitutions_fa
	'it': substitutions_it
	'nl': substitutions_nl
	'no': substitutions_no
	'ru': substitutions_ru
}
