module slugify

const substitutions_ru = {
	'а':  'a'
	'б':  'b'
	'в':  'v'
	'г':  'g'
	'д':  'd'
	'е':  'e'
	'ё':  'yo'
	'ж':  'zh'
	'з':  'z'
	'дж': 'j'
	'и':  'i'
	'й':  'y'
	'к':  'k'
	'л':  'l'
	'м':  'm'
	'н':  'n'
	'о':  'o'
	'п':  'p'
	'р':  'r'
	'с':  's'
	'т':  't'
	'у':  'u'
	'ф':  'f'
	'х':  'h'
	'ц':  'ts'
	'ч':  'ch'
	'ш':  'sh'
	'щ':  'sch'
	'ъ':  ''
	'ы':  'i'
	'ь':  ''
	'э':  'e'
	'ю':  'yu'
	'я':  'ya'
	'%':  'procent'
	'♥':  'serdtse'
	'&':  'i'
	'@':  'sobaka'
	'#':  'reshyotka'
	'=':  'ravno'
	'~':  'tilda'
	'<':  'menshe'
	'>':  'bolshe'
	'|':  'ili'
	'∞':  'beskonechnost'
}
