module slugify

const substitutions_fa = {
	'ک': 'kh'
	'ی': 'y'
}
