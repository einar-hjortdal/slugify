module slugify

const substitutions_nl = {
	'&': 'en'
	'@': 'at'
}
