module slugify

const substitutions_it = {
	'&': 'e'
	'@': 'chiocciola'
	'%': 'per cento'
	'<': 'minore'
	'>': 'maggiore'
	'|': 'o'
}
